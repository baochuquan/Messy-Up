module test;
wire C;
wire [3:0] sum;
reg [3:0] X;
reg [3:0] Y;

add_4 hhd(.X(X), .Y(Y), .sum(sum), .C(C));
initial begin
		
end
endmodule
